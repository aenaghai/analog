magic
tech scmos
timestamp 1668061076
<< error_p >>
rect -21 15 31 16
rect -22 12 -21 15
rect -7 12 1 15
rect 3 12 10 15
rect 11 12 15 15
rect 31 12 32 15
rect -21 11 -7 12
rect -5 11 -3 12
rect -1 11 3 12
rect 5 11 6 12
rect 8 11 11 12
rect 13 11 31 12
rect -8 9 -4 11
rect -1 10 1 11
rect 10 9 12 10
rect -21 8 22 9
rect -6 7 -3 8
rect 10 7 12 8
rect -1 6 0 7
rect 12 6 14 7
rect -3 5 0 6
rect -4 3 -3 5
rect -1 4 3 5
rect 9 4 10 6
rect 12 4 13 6
rect -1 3 4 4
rect -3 2 0 3
rect 2 2 4 3
rect 9 2 13 4
rect -21 1 22 2
rect -2 0 0 1
rect 12 0 14 1
rect 0 -1 2 0
rect 3 -1 4 0
rect -3 -15 -2 -1
rect 0 -14 1 -1
rect 3 -2 6 -1
rect 3 -3 7 -2
rect 4 -4 7 -3
rect 4 -5 6 -4
rect 0 -15 3 -14
rect -3 -16 1 -15
rect 5 -16 7 -15
rect -3 -17 7 -16
rect -3 -18 -2 -17
rect 0 -18 2 -17
rect -3 -19 2 -18
rect 5 -19 6 -18
rect 1 -20 3 -19
rect -1 -21 3 -20
rect 4 -21 6 -19
rect -2 -22 -1 -21
rect 1 -22 6 -21
rect -2 -23 6 -22
rect -1 -25 3 -23
rect 4 -25 6 -23
rect -2 -26 6 -25
rect 7 -19 9 -17
rect 7 -26 8 -19
rect -2 -28 8 -26
rect -3 -37 -2 -28
rect 0 -30 2 -28
rect 7 -30 9 -28
rect 0 -37 1 -30
rect -13 -38 -11 -37
rect -3 -38 1 -37
rect 3 -38 5 -37
rect 11 -38 13 -37
rect -22 -39 31 -38
rect -23 -41 -22 -39
rect -13 -41 -9 -39
rect -2 -41 2 -39
rect 3 -41 7 -39
rect 11 -41 15 -39
rect 31 -41 32 -39
rect -22 -42 -13 -41
rect -11 -42 -2 -41
rect 0 -42 3 -41
rect 5 -42 11 -41
rect 13 -42 31 -41
<< nwell >>
rect -27 -10 35 29
<< ntransistor >>
rect 1 -19 3 -17
rect 1 -30 3 -28
<< ptransistor >>
rect -1 6 1 8
rect 2 -1 4 1
<< ndiffusion >>
rect 0 -19 1 -17
rect 3 -19 5 -17
rect 0 -30 1 -28
rect 3 -30 5 -28
<< pdiffusion >>
rect -21 7 -7 8
rect -5 7 -1 8
rect -21 6 -1 7
rect 1 7 22 8
rect 1 6 10 7
rect 12 6 22 7
rect -21 0 2 1
rect -21 -1 -2 0
rect 0 -1 2 0
rect 4 0 10 1
rect 12 0 22 1
rect 4 -1 22 0
<< ndcontact >>
rect -2 -19 0 -17
rect 5 -19 7 -17
rect -2 -30 0 -28
rect 5 -30 7 -28
<< pdcontact >>
rect -7 7 -5 8
rect 10 6 12 7
rect -2 -1 0 0
rect 10 0 12 1
<< psubstratepcontact >>
rect -13 -41 -11 -39
rect -2 -41 0 -39
rect 3 -41 5 -39
rect 11 -41 13 -39
<< nsubstratencontact >>
rect -7 12 -5 15
rect -3 12 -1 15
rect 3 12 5 15
rect 6 12 8 15
rect 11 12 13 15
<< polysilicon >>
rect -1 8 1 10
rect -1 5 1 6
rect 0 3 1 5
rect 2 1 4 2
rect 2 -2 4 -1
rect 2 -4 3 -2
rect 1 -17 3 -15
rect 1 -21 3 -19
rect 1 -28 3 -27
rect 1 -33 3 -30
<< polycontact >>
rect -1 3 0 5
rect 3 -4 4 -2
rect 1 -23 3 -21
rect 1 -27 3 -25
<< rmetal1 >>
rect -21 12 -7 15
rect -5 12 -3 15
rect -1 12 3 15
rect 5 12 6 15
rect 8 12 11 15
rect 13 12 31 15
rect -7 8 -5 12
rect -3 3 -1 5
rect 10 1 12 6
rect -2 -17 0 -1
rect 4 -4 6 -2
rect -1 -23 1 -21
rect -1 -27 1 -25
rect 5 -28 7 -19
rect -2 -39 0 -30
rect -22 -41 -13 -39
rect -11 -41 -2 -39
rect 0 -41 3 -39
rect 5 -41 11 -39
rect 13 -41 31 -39
<< labels >>
rlabel rmetal1 -11 14 -11 14 1 Vdd
rlabel rmetal1 -18 -40 -18 -40 1 gnd
rlabel rmetal1 -2 4 -2 4 1 Vbias1
rlabel rmetal1 5 -3 5 -3 1 Vbias2
rlabel rmetal1 0 -22 0 -22 1 Vbias3
rlabel rmetal1 0 -26 0 -26 1 Vs
rlabel rmetal1 -1 -12 -1 -12 1 Vout
<< end >>
